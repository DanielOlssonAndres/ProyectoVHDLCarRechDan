library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity TOP_tb is
end TOP_tb;


architecture Behavioral of TOP_tb is
begin

end architecture;
