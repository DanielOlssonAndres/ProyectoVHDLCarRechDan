library ieee;
use ieee.std_logic_1164.ALL;

entity decod_display_tb is
end decod_display_tb;

architecture Behavioral of decod_display_tb is

begin


end Behavioral;
