library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--use IEEE.NUMERIC_STD.ALL;

entity Controlador_de_Sec_tb is
end entity;

architecture Behavioral of Controlador_de_Sec is

begin

end architecture;