library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity TOP is

end TOP;

architecture STRUCTURAL of TOP is

begin

end architecture;
