library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package paquete_types is
    type vec_integrer is array(natural range <>) of integer;
end paquete_types;
